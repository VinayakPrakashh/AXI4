module APB_MASTER #(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 32
) (
    input PCLK,
    input PRESETn,
    // APB Master Interface
    output reg PSEL_UART,
    output reg PSEL_TIMER,
    output reg PENABLE,
    output reg PWRITE,
    output reg [ADDR_WIDTH-1:0] PADDR,
    output reg [DATA_WIDTH-1:0] PWDATA,
    input [DATA_WIDTH-1:0] PRDATA,
    input PREADY,
    input PSLVERR,
    // Control signals AXI4 to APB
    input transfer,
    input read,
    input write,
    // axi4 inputs for simulation purposes
    input [ADDR_WIDTH-1:0] apb_waddr,
    input [ADDR_WIDTH-1:0] apb_raddr,
    input [DATA_WIDTH-1:0] apb_wdata,
    output reg [DATA_WIDTH-1:0] apb_rdata
);

wire error;
reg [1:0] state, next_state;

parameter IDLE = 2'b00,
          SETUP = 2'b01,
          ACCESS = 2'b10;
always @(posedge PCLK) begin
    if (!PRESETn)
        state <= IDLE;
    else
        state <= next_state; 
end

always @(*) begin
    case (state)
    IDLE: begin
        if (transfer) // Start condition
            next_state = SETUP;
        else
            next_state = IDLE;
    end
    SETUP:
        next_state = ACCESS;
    ACCESS: begin
        if (PREADY && !transfer)
            next_state = IDLE;
        else if(PREADY && transfer)
            next_state = SETUP;
        else
            next_state = ACCESS;
    end
    endcase
end

always @(state) begin
 case (state)
    IDLE: begin
        PSEL_UART <= 1'b0;
        PSEL_TIMER <= 1'b0;
        PENABLE <= 1'b0;
    end 
    SETUP: begin
        PSEL_UART <= (apb_waddr[ADDR_WIDTH-1:ADDR_WIDTH-4] == 0) ? 1'b1 : 1'b0;
        PSEL_TIMER <= (apb_waddr[ADDR_WIDTH-1:ADDR_WIDTH-4] > 0) ? 1'b1 : 1'b0;
        PENABLE <= 1'b0;
        if(write) begin
            PWRITE <= 1'b1;
            PADDR <= apb_waddr;
            PWDATA <= apb_wdata;
        end else if(read) begin
            PWRITE <= 1'b0;
            PADDR <= apb_raddr;
        end
    end
    ACCESS: begin
        PENABLE <= 1'b1;
        if(!PWRITE && PREADY) begin
            apb_rdata <= PRDATA;
        end
    end
    default: begin
        PSEL_UART <= 1'b0;
        PSEL_TIMER <= 1'b0;
        PENABLE <= 1'b0;
    end
 endcase
    end


assign error = PSLVERR & (PSEL_UART | PSEL_TIMER) & PENABLE; //just for future use
endmodule